module fourbitadder (input logic [3:0], output logic [4:0] sum);


endmodule