module fourbitadder (input logic [3:0] a, input logic [3:0] b, output logic [4:0] sum);
	assign sum = a + b;
	
//	logic [3:0] c;
//	always_comb
//		sum[0] <= a[0] ^ b[0];
//		c[0] <= a[0] & b[0];
		
//		sum[1] <= (a[1] ^ b[1]) ^ c[0];
//		c[1] <= (a[1] & b[1]) | (a[1] & c[0]) | (b[1] & c[0]);
		
		
//		sum[2] <= (a[2] ^ b[2]) ^ c[1];
//		c[2] <= (a[2] & b[2]) | (a[2] & c[1]) | (b[2] & c[1]);
		
//		
//		sum[3] <= (a[3] ^ b[3]) ^ c[1];
//		c[3] <= (a[3] & b[3]) | (a[3] & c[3]) | (b[3] & c[2]);
		
		
//		sum[4] <= (a[4] ^ b[4]) ^ c[3];
//		c[4] <= (a[4] & b[4]) | (a[4] & c[4]) | (b[4] & c[3]);
		
		
//		sum[5] <= c[4];
	
endmodule
