module keypad_getrowcol(
	input logic [31:0] counter; // what frequency to write row high and read col, then switch
	input logic [3:0] rows;
	output logic [3:0] cols;
);





endmodule